* DIODE COMPARISON
* Second Input Deck

VDD VIN 0
D1 VIN 0 D1
D2 VIN 0 D2
D3 VIN 0 D3


.MODEL D1 D RS=1 IS=1E-14
.MODEL D2 D RS=1 IS=1E-13
.MODEL D3 D RS=1 IS=1E-12

.DC VDD 0 2 0.01

.PROBE
.PRINT DC I(D1) I(D2) I(D3)
.END
